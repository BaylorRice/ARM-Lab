`timescale 1ns / 1ps
`include "definitions.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 02/12/2024 01:50:24 PM
// Design Name: Register File
// Module Name: regfile
// Project Name: Lab 4 - Beginnning to Decode
// Target Devices: Vivado Simulation
// Tool Versions: Vivado 2021.2
// Description: *shrug*
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module regfile(

    );
endmodule
