`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 03/25/2024 12:28:52 PM
// Design Name: Aritmatic Logic Unit ("ALU")
// Module Name: alu
// Project Name: Lab 8 - ALU and ALU Control
// Target Devices: Vivado Simulator
// Tool Versions: Vivado 2021.2
// Description: figure it out
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module alu(

    );
endmodule
