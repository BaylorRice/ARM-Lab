`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 02/19/2024 12:30:48 PM
// Design Name: Control Unit
// Module Name: control
// Project Name: Lab 5 - Control Unit and Sign Extender
// Target Devices: Vivado Simulation
// Tool Versions: Vivado 2021.2
// Description: Who cares
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control(

    );
endmodule
