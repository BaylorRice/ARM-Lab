`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 02/19/2024 01:47:03 PM
// Design Name: Sign Extender
// Module Name: sign_extender
// Project Name: Lab 5 - Control unit and Sign Extenders
// Target Devices: Vivado Simulation
// Tool Versions: Vivado 2021.2
// Description: figure it out
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module sign_extender(
    input [`INSTR_LEN-1:0] instruction,
    output reg [`WORD-1:0] sign_extended_output
    );
    
    
endmodule
