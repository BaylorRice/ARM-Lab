`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 02/26/2024 12:34:43 PM
// Design Name: Decode Stage Wrapper Module
// Module Name: iDecode
// Project Name: Lab 6 - Finishing Decode
// Target Devices: Vivado Simulation
// Tool Versions: Vivado 2021.2
// Description: See Pg. 28 of the manual, I mean, figure it out.
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module iDecode(
    input wire
    );
endmodule
