`timescale 1ns / 1ps
`include "definitions.vh"
//////////////////////////////////////////////////////////////////////////////////
// Company: Baylor University
// Engineer: Reese Ford
// 
// Create Date: 03/28/2024 12:55:30 PM
// Design Name: Instruction Execution Wrapper
// Module Name: iExecute
// Project Name: Lab 9 - Execute Stage
// Target Devices: Vivado Simulator
// Tool Versions: Vivado 2021.2
// Description: beats me
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module iExecute(

    );
endmodule
